`include "risc_v_pipeline_define.svh"
module control (
    input            clk            ,
    input            rst_n          ,
    input            BrEq_i         ,
    input            BrLT_i         ,
    input      [6:0] opcode_i       ,
    input      [6:0] funct7_i       ,
    input      [2:0] funct3_i       ,
    output reg [2:0] ImmSel_o       ,
    output reg       PCSel_o        ,
    output reg       BrUn_o         ,
    output reg       ASel_o         ,
    output reg       BSel_o         ,
    output reg       MemRW_o        ,
    output reg       RegWEn_o       ,
    output reg [1:0] WBSel_o        ,
    output reg [3:0] ALUSel_o       ,
    output           insert_nop_flag
);
  reg PCSel;

  //insert 2 nop for JAL
  reg  count          ;
  wire detect_jal     ;
  wire pc_sel_jal     ;
  reg  pc_sel_jal_reg ;

  assign detect_jal = (opcode_i == `J);

  always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
      count <= 0;
    end else if(detect_jal) begin
      count <= count + 1;
    end else begin
      count <= 0;
    end
  end

  assign insert_nop_flag = detect_jal || (count == 1'b1);

  always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
      pc_sel_jal_reg <= 0;
    end else begin
      pc_sel_jal_reg <= pc_sel_jal;
    end
  end

  assign PCSel_o = (count == 1) ? pc_sel_jal_reg : PCSel;

  // Control logic
  always @(*)
  begin
      case(opcode_i)
      `R:
          case(funct3_i)
          3'b000:
              case(funct7_i)
              7'b0000000: //add
                  begin
                      PCSel       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      //BrUn_o        = 1'b0;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUadd;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              7'b0100000: //sub
                  begin
                      PCSel       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      //BrUn_o        = 1'b0;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsub;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              endcase
          3'b001: //sll
              begin
                  PCSel           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUsll;
                  MemRW_o           = 0;//Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b010: //slt
              begin
                  PCSel           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUslt;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b011: //sltu
              begin
                  PCSel           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUsltu;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b100: //xor
              begin
                  PCSel           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUxor;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b101:
              case(funct7_i)
              7'b0000000: //srl
                  begin
                      PCSel       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      // BrUn_o        = 1'bx;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsrl;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              7'b0100000: //sra
                  begin
                      PCSel       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      // BrUn_o        = 1'bx;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsra;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              endcase
          3'b110: //or
              begin
                  PCSel           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUor;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b111: //and
              begin
                  PCSel           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUand;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          endcase
      `IMM_I:
        begin
            PCSel               = 0; //PC=PC+4
            ImmSel              = ImmSelI; //Immediate type I
            // BrUn                = 1'bx;
            ASel                = 0; //Reg
            BSel                = 1; //Imm
            ALUSel              = ALUadd;
            MemRW               = 0; //Read
            RegWEn              = 1;
            WBSel               = 2'b01; //ALU
        end
      `LOAD_I:
          begin
              PCSel               = 0; //PC=PC+4
              ImmSel_o              = `ImmSelI; //Immediate type I
              BrUn_o                = 1'bx;
              ASel_o                = 0; //Reg
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b00; //Mem
              end
      `S:
          begin
              PCSel               = 0; //PC=PC+4
              ImmSel_o              = `ImmSelS; //Immediate type S
              BrUn_o                = 1'bx;
              ASel_o                = 0; //Reg
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 1; //Write
              RegWEn_o              = 0;
              WBSel_o               = 2'bxx;
              end
      `B:
          case(funct3_i)
          3'b000: //beq // Branchcomp block read BrEq_i and change PCSel
              begin
                  PCSel           = (BrEq_i) ? 1 : 0; //PC=PC+Imm when Eq, PC= PC+4 when not Eq
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  // BrUn_o            = 1'bx;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          3'b001: //bne //Branchcomp read BrEq_i and change PCSel
              begin
                  PCSel           = (BrLT_i) ? 0 : 1; //ALU // temporary value
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  // BrUn_o            = 1'bx;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          3'b100: //blt //Branchcomp read BrLT_i and change PCSel
              begin
                  PCSel           = (BrLT_i) ? 1 : 0; //PC+4 // temporary value
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  BrUn_o            = 0;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0;//Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          3'b101: //bltu //Branchcomp read BrLT_i and change PCSel
              begin
                  PCSel           = (BrLT_i) ? 1 : 0; //PC+4 // temporary value
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  BrUn_o            = 1;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          endcase
      `JUMP_I:
          begin
              PCSel               = 2; //jump_pc
              ImmSel_o              = `ImmSelI; //Immediate type I
              // BrUn_o                = 1'bx;
              ASel_o                = 0; //Reg
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b10; // PC+4
          end
      `J:
          begin
              pc_sel_jal            = 1; //jump_pc
              ImmSel_o              = `ImmSelJ; //Immediate type J
              ASel_o                = 1; //PC
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b10; // PC+4
          end
      `U:
          begin
              PCSel               = 0; //PC+4
              ImmSel_o              = `ImmSelU; //Immediate type U
              BrUn_o                = 1'bx;
              ASel_o                = 1; //PC
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b01; // ALU
          end

      default: 
        begin
              PCSel                 = 0; //PC+4
              ImmSel_o              = 4'b1111;
              BrUn_o                = 0;
              ASel_o                = 0; //PC
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUnop;
              MemRW_o               = 0; //Read
              RegWEn_o              = 0;
              WBSel_o               = 2'b01; // ALU
        end
      endcase
  end
endmodule
