module risc_v_pipeline (
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	
);

endmodule : risc_v_pipeline