`include "risc_v_pipeline_define.svh"
module control (
    input            clk      ,
    input            rst_n    ,
    input            BrEq_i   ,
    input            BrLT_i   ,
    input      [6:0] opcode_i ,
    input      [6:0] funct7_i ,
    input      [2:0] funct3_i ,
    output reg [2:0] ImmSel_o ,
    output reg       PCSel_o  ,
    output reg       BrUn_o   ,
    output reg       ASel_o   ,
    output reg       BSel_o   ,
    output reg       MemRW_o  ,
    output reg       RegWEn_o ,
    output reg [1:0] WBSel_o  ,
    output reg [3:0] ALUSel_o  
);

  always @(*)
  begin
      case(opcode_i)
      `R:
          case(funct3_i)
          3'b000:
              case(funct7_i)
              7'b0000000: //add
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      //BrUn_o        = 1'b0;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUadd;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              7'b0100000: //sub
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      //BrUn_o        = 1'b0;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsub;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              endcase
          3'b001: //sll
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUsll;
                  MemRW_o           = 0;//Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b010: //slt
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUslt;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b011: //sltu
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUsltu;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b100: //xor
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUxor;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b101:
              case(funct7_i)
              7'b0000000: //srl
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      // BrUn_o        = 1'bx;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsrl;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              7'b0100000: //sra
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      // BrUn_o        = 1'bx;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsra;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              endcase
          3'b110: //or
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUor;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b111: //and
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUand;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          endcase
      `IMM_I:
          case(funct3_i)
          3'b000:
              case(funct7_i)
              7'b0000000: //add
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      //BrUn_o        = 1'b0;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUadd;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              7'b0100000: //sub
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      //BrUn_o        = 1'b0;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsub;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              endcase
          3'b001: //sll
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUsll;
                  MemRW_o           = 0;//Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b010: //slt
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUslt;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b011: //sltu
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUsltu;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b100: //xor
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUxor;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b101:
              case(funct7_i)
              7'b0000000: //srl
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      // BrUn_o        = 1'bx;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsrl;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              7'b0100000: //sra
                  begin
                      PCSel_o       = 0; //PC=PC+4
                      ImmSel_o      = `ImmSelR;
                      // BrUn_o        = 1'bx;
                      ASel_o        = 0; //Reg
                      BSel_o        = 0; //Reg
                      ALUSel_o      = `ALUsra;
                      MemRW_o       = 0; //Read
                      RegWEn_o      = 1;
                      WBSel_o       = 2'b01; //ALU
                  end
              endcase
          3'b110: //or
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUor;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          3'b111: //and
              begin
                  PCSel_o           = 0; //PC=PC+4
                  ImmSel_o          = `ImmSelR;
                  // BrUn_o            = 1'bx;
                  ASel_o            = 0; //Reg
                  BSel_o            = 0; //Reg
                  ALUSel_o          = `ALUand;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 1;
                  WBSel_o           = 2'b01; //ALU
              end
          endcase
      `LOAD_I:
          begin
              PCSel_o               = 0; //PC=PC+4
              ImmSel_o              = `ImmSelI; //Immediate type I
              BrUn_o                = 1'bx;
              ASel_o                = 0; //Reg
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b00; //Mem
              end
      `S:
          begin
              PCSel_o               = 0; //PC=PC+4
              ImmSel_o              = `ImmSelS; //Immediate type S
              BrUn_o                = 1'bx;
              ASel_o                = 0; //Reg
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 1; //Write
              RegWEn_o              = 0;
              WBSel_o               = 2'bxx;
              end
      `B:
          case(funct3_i)
          3'b000: //beq // Branchcomp block read BrEq_i and change PCSel_o
              begin
                  PCSel_o           = (BrEq_i) ? 1 : 0; //PC=PC+Imm when Eq, PC= PC+4 when not Eq
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  // BrUn_o            = 1'bx;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          3'b001: //bne //Branchcomp read BrEq_i and change PCSel_o
              begin
                  PCSel_o           = (BrLT_i) ? 0 : 1; //ALU // temporary value
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  // BrUn_o            = 1'bx;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          3'b100: //blt //Branchcomp read BrLT_i and change PCSel_o
              begin
                  PCSel_o           = (BrLT_i) ? 1 : 0; //PC+4 // temporary value
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  BrUn_o            = 0;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0;//Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          3'b101: //bltu //Branchcomp read BrLT_i and change PCSel_o
              begin
                  PCSel_o           = (BrLT_i) ? 1 : 0; //PC+4 // temporary value
                  ImmSel_o          = `ImmSelB; //Immediate type `B
                  BrUn_o            = 1;
                  ASel_o            = 1; //PC
                  BSel_o            = 1; //Imm
                  ALUSel_o          = `ALUadd;
                  MemRW_o           = 0; //Read
                  RegWEn_o          = 0;
                  WBSel_o           = 2'bxx;
              end
          endcase
      `JUMP_I:
          begin
              PCSel_o               = 2; //jump_pc
              ImmSel_o              = `ImmSelI; //Immediate type I
              // BrUn_o                = 1'bx;
              ASel_o                = 0; //Reg
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b10; // PC+4
          end
      `J:
          begin
              PCSel_o               = 1; //jump_pc
              ImmSel_o              = `ImmSelJ; //Immediate type J
              ASel_o                = 1; //PC
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b10; // PC+4
          end
      `U:
          begin
              PCSel_o               = 0; //PC+4
              ImmSel_o              = `ImmSelU; //Immediate type U
              BrUn_o                = 1'bx;
              ASel_o                = 1; //PC
              BSel_o                = 1; //Imm
              ALUSel_o              = `ALUadd;
              MemRW_o               = 0; //Read
              RegWEn_o              = 1;
              WBSel_o               = 2'b01; // ALU
          end

      default: ALUSel_o             = `ALUnop;
      endcase
  end
endmodule
